module four_bit_adder_testbench;

	reg [3:0] a;
	reg [3:0] b;
	wire [3:0] sum;
     wire finalcarry;

	four_bit_adder testbench (
  	  .a(a),
  	  .b(b),
  	  .sum(sum),
   	  .finalcarry(finalcarry)
	);
    
	integer i,j,k;
   // $dumpfile("dump.vcd"); $dumpvars;
	initial begin
  	  $display("a    b   finalcarry    sum");
      $monitor("%b %b %b %b %b", a, b, finalcarry, sum);
   		 for (i = 0; i < 16; i = i + 1) begin
   			 for (j = 0; j < 16; j = j + 1) begin
   				  a=i;
  				  b=j;
  				  #10;
   			 end
   		 end
  	  $finish;
    end

endmodule
