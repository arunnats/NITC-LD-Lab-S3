module fourBitDecrementor(
	input [3:0] a,
	output [4:0] b
);
    wire [3:0]carry;
    
    fullAdder fa0(.s(b[0]),.c(carry[0]),.a(a[0]),.b(1'b1),.cin(1'b0));
    fullAdder fa1(.s(b[1]),.c(carry[1]),.a(a[1]),.b(1'b1),.cin(carry[0]));
    fullAdder fa2(.s(b[2]),.c(carry[2]),.a(a[2]),.b(1'b1),.cin(carry[1]));
    fullAdder fa3(.s(b[3]),.c(carry[3]),.a(a[3]),.b(1'b1),.cin(carry[2]));
    
    not_1In not_1 (b[4],carry[3]);
    
endmodule

module and_2In(
	output y,
	input a,
   b
);
    
	wire aNandb;
    
	nand nand_1 (aNandb,a,b);
	nand nand_2 (y,aNandb,aNandb);

endmodule

module or_2In(
	output y,
	input a,
	input b
);
    
	wire aNanda, bNandb;
    
	nand nand_1 (aNanda,a,a);
	nand nand_2 (bNandb,b,b);
	nand nand_3 (y,aNanda,bNandb);

endmodule

module not_1In(
	output y,
	input a
);
    
	nand nand_1 (y,a);
    
endmodule

module xor_2In(
	output y,
	input a,
	b
);

	wire aNandb,aNandComp,bNandComp;

	nand nand_1 (aNandb,a,b);
	nand nand_2 (aNandComp,a,aNandb);
	nand nand_3 (bNandComp,b,aNandb);
	nand nand_4 (y,aNandComp,bNandComp);

endmodule

module halfAdder(
	output s,
	c,
	input a,
	b
);

	xor_2In xor_1(.y(s),.a(a),.b(b));
	and_2In and_1(.y(c),.a(a),.b(b));
    
endmodule

module fullAdder(
    output s,
    c,
    input a,
    b,
    cin
);
    
    wire carry1,carry2,sum;
    halfAdder ha1(.s(sum),.c(carry1),.a(a),.b(b));
    halfAdder ha2(.s(s),.c(carry2),.a(cin),.b(sum));
    
    or_2In or1(c,carry1,carry2);
    
endmodule
