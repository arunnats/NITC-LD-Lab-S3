module bcd_adder_test();
	 reg [3:0] a,
    reg [3:0] b,
    wire [3:0] sum,
    wire finalcarry
	 
	 bcd_adder testbench(
  	  .a(a),
  	  .b(b),
  	  .sum(sum),
     .finalcarry(finalcarry)
	);
	
	integer i,j;
    
	initial begin
  	  $display("a    b	finalcarry    sum");
  	  $monitor("%b %b %b %b", a, b, finalcarry, sum);
   	  for (k = 0; k < 9; k = k + 1) begin
   		 for (i = 0; i < 9; i = i + 1) begin
   			  a=i;
  				  b=j;
  				  #10;
   		 end
   	 end
  	  $finish;
    end
endmodule
