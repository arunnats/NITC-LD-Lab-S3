module bcd_excess3_test();
  reg [3:0]a;
  wire [3:0]e;
  
  bcd_excess3 uut (.a(a),.e(e));
 
  integer count;
  
  initial begin
    for(count=0;count<16;count=count+1) begin
      {a}=count;
      #10;
    end
	 end
	 endmodule