module bcd_adder_testbench;

   reg [3:0] a;
   reg [3:0] b;
   wire [3:0] sum;
   wire finalcarry;

   bcd_adder testbench (
    	.a(a),
    	.b(b),
    	.sum(sum),
    .   	 finalcarry(finalcarry));
    
	integer i,j;
    
	initial begin
	//$display("a    b    finalcarry    sum");
    //	$monitor("%b %b %b %b", a, b, finalcarry, sum);
     	   for (i = 0; i < 10; i = i + 1) begin
     		   for (j = 0; j < 10; j = j + 1) begin
     				a=i;
				  	 b=j;
					#10;
     		   end
     	   end

    	$finish;
    end

endmodule
